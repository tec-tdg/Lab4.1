module Sumador_punto_flotante_tb();




endmodule 